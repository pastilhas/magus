module main

import www

fn main() {
	www.run()
}
