module main

struct Author {
	name string
}
