module main

struct Tag {
	name string
}
