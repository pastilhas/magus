module main

fn main() {
	run()
}
